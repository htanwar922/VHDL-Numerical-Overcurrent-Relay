
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use std.textio.all;
use ieee.std_logic_textio.all;

use work.my_functions.all;
use work.my_types.all;

package my_fixed_package is



end my_fixed_package;


package body my_fixed_package is



end my_fixed_package;