
library ieee;
use ieee.std_logic_1164.all;
use std.textio.all;

use work.my_types.all;
use work.my_float_package.all;
use work.my_functions.all;

entity dft32 is
	generic( N : natural := 40 );
	port (
        clk : in std_logic := '0';
        adc : in float32;
        X_1 : out float32
    );
end entity;

architecture dft32 of dft32 is
	signal C : float32_arr(0 to N-1+N/4) :=
		(
				"00000000000000000000000000000000",
            "00111110001000000011000001011000",
            "00111110100111100011011101111000",
            "00111110111010000111000101110000",
            "00111111000101100111100100011000",
            "00111111001101010000010011110010",
            "00111111010011110001101110111100",
            "00111111011001000001100100000000",
            "00111111011100110111100001110000",
            "00111111011111001101100100100100",
            "00111111100000000000000000000000",
            "00111111011111001101100100100100",
            "00111111011100110111100001110000",
            "00111111011001000001100100000000",
            "00111111010011110001101110111100",
            "00111111001101010000010011110010",
            "00111111000101100111100100011000",
            "00111110111010000111000101110000",
            "00111110100111100011011101111000",
            "00111110001000000011000001011000",
            "00000000000000000000000000000000",
            "10111110001000000011000001011000",
            "10111110100111100011011101111000",
            "10111110111010000111000101110000",
            "10111111000101100111100100011000",
            "10111111001101010000010011110010",
            "10111111010011110001101110111100",
            "10111111011001000001100100000000",
            "10111111011100110111100001110000",
            "10111111011111001101100100100100",
            "10111111100000000000000000000000",
            "10111111011111001101100100100100",
            "10111111011100110111100001110000",
            "10111111011001000001100100000000",
            "10111111010011110001101110111100",
            "10111111001101010000010011110010",
            "10111111000101100111100100011000",
            "10111110111010000111000101110000",
            "10111110100111100011011101111000",
            "10111110001000000011000001011000",
            "00000000000000000000000000000000",
            "00111110001000000011000001011000",
            "00111110100111100011011101111000",
            "00111110111010000111000101110000",
            "00111111000101100111100100011000",
            "00111111001101010000010011110010",
            "00111111010011110001101110111100",
            "00111111011001000001100100000000",
            "00111111011100110111100001110000",
            "00111111011111001101100100100100"
		);
	signal N_float     : float32 := b"0_1000_0100_0100_0000_0000_0000_0000_000";
	signal two_float   : float32 := b"0_1000_0000_0000_0000_0000_0000_0000_000";
	signal x   : float32_arr(0 to N-1);
	signal tmp 	: float32 := b"0_0111_1111_0000_0000_0000_0000_0000_000";
begin
	
	process_calculate_X1 : process(clk)
        variable tmp_S 	: float32 := b"0_0000_0000_0000_0000_0000_0000_0000_000";
        variable tmp_C 	: float32 := b"0_0000_0000_0000_0000_0000_0000_0000_000";
        variable sqrt_tmp 	: float32 := b"0_0111_1111_0000_0000_0000_0000_0000_000";
	begin
		if rising_edge(clk) then
			for i in 0 to N-1 loop
				tmp_S := tmp_S + x(i) * C(i);
				tmp_C := tmp_C + x(i) * C(i + N/4);
			end loop;
		end if;
		if falling_edge(clk) then
            tmp <= tmp_S * two_float;
		end if;
		X_1 <= sqrt(tmp);
	end process;
	
--	process_update_samples : process(clk, x)
--        variable current : natural := 0;
--	begin
----		if rising_edge(clk) then
----			x(current) <= adc;
----			current := current+1;
----			if(current = N) then current := 0; end if;
----		end if;
--	end process;
	
end architecture;